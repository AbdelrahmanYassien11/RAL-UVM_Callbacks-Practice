package pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
  
    `include "seq_item.sv"
    `include "ral_pkg.sv"
    `include "ral2axi_adapter.sv"

    `include "base_seq.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "agent.sv"
    `include "env.sv"
    `include "base_test.sv"
endpackage : pkg